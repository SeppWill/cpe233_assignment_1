module cntr_udclr_nb(clk, clr, up, ld, D, count, rco);
	input   clk, clr, up, ld;
	input   [n-1:0] D;
	output  reg [n-1:0] count;
	output  reg rco;

	//- default data-width

	parameter n = 8;

	always @(posedge clr, posedge clk)
	begin
		if (clr == 1)       // asynch reset count <= 0;
		else if (ld == 1)   // load new value count <= D;
		else if (up == 1)   // count up (increment) count <= count + 1;
		else if (up == 0)   // count down (decrement) count <= count - 1;
	end

	//- handles the RCO, which is direction dependent

	always @(count, up)
	begin
		if ( up == 1 && &count == 1'b1) rco = 1'b1;
		else if (up == 0 && |count == 1'b1) rco = 1'b1;
		else
			rco = 1'b0;

	end
endmodule


